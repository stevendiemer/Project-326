`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:10:59 03/08/2012 
// Design Name: 
// Module Name:    game_message 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module game_message(
    input [3:0] coins_left,
	 input [10:0] hcount, 
	 input [10:0] vcount,
	 input clk,
	 input rst,
    output r,
    output g,
    output b
    );


endmodule
