`timescale 1ns / 1ps
// ------------------------------------------------------------------------
// vga_controller_640_60.vhd
//----------------------------------------------------------------------
// Author : Chirag Parikh
//          
//----------------------------------------------------------------------
// Software version : Xilinx ISE 10.1.03i
//                    WebPack
// Device	        : xc3s500e-4fg320
// ------------------------------------------------------------------------
// This file contains the logic to generate the synchronization signals,
// horizontal and vertical pixel counter and video disable signal
// for the 640x480@60Hz resolution.
// ------------------------------------------------------------------------
//  Behavioral description
// ------------------------------------------------------------------------
// Please read the following article on the web regarding the vga video timings:
// http://www.epanorama.net/documents/pc/vga_timing.html

// This module generates the video synch pulses for the monitor to
// enter 640x480@60Hz resolution state. It also provides horizontal
// and vertical counters for the currently displayed pixel and a blank
// signal that is active when the pixel is not inside the visible screen
// and the color outputs should be reset to 0.

// timing diagram for the horizontal synch signal (HS)
// 0                         648    744           800 (pixels)
// -------------------------|______|-----------------
// timing diagram for the vertical synch signal (VS)
// 0                                  482    484  525 (lines)
// -----------------------------------|______|-------

// The blank signal is delayed one pixel clock period (40ns) from where
// the pixel leaves the visible screen, according to the counters, to
// account for the pixel pipeline delay. This delay happens because
// it takes time from when the counters indicate current pixel should
// be displayed to when the color data actually arrives at the monitor
// pins (memory read delays, synchronization delays).
// ------------------------------------------------------------------------
//  Port definitions
// ------------------------------------------------------------------------
// rst               - global reset signal
// pixel_clk         - input pin, from dcm_25MHz
//                   - the clock signal generated by a DCM that has
//                   - a frequency of 25MHz.
// HS                - output pin, to monitor
//                   - horizontal synch pulse
// VS                - output pin, to monitor
//                   - vertical synch pulse
// hcount            - output pin, 11 bits, to clients
//                   - horizontal count of the currently displayed
//                   - pixel (even if not in visible area)
// vcount            - output pin, 11 bits, to clients
//                   - vertical count of the currently active video
//                   - line (even if not in visible area)
// blank             - output pin, to clients
//                   - active when pixel is not in visible area.
// ------------------------------------------------------------------------


// the vga_controller_640_60 module declaration
// read above for behavioral description and port definitions.
module vga_controller_640_60(rst, pixel_clk, HS, VS, hcount, vcount, blank);

input rst, pixel_clk;
output HS, VS;
output [10:0]hcount, vcount;
output blank;

// ------------------------------------------------------------------------
// CONSTANTS
// ------------------------------------------------------------------------

// maximum value for the horizontal pixel counter
parameter HMAX = 11'b01100100000;                             // 800
// maximum value for the vertical pixel counter
parameter VMAX = 11'b01000001101;                             // 525
// total number of visible columns
parameter HLINES = 11'b01010000000;                           // 640
// value for the horizontal counter where front porch ends
parameter HFP = 11'b01010001000;                              // 648
// value for the horizontal counter where the synch pulse ends
parameter HSP = 11'b01011101000;                              // 744
// total number of visible lines
parameter VLINES = 11'b00111100000;                           // 480
// value for the vertical counter where the front porch ends
parameter VFP = 11'b00111100010;                              // 482
// value for the vertical counter where the synch pulse ends
parameter VSP = 11'b00111100100;                              // 484
// polarity of the horizontal and vertical synch pulse
// only one polarity used, because for this resolution they coincide.
parameter SPP = 1'b0;


// ------------------------------------------------------------------------
// SIGNALS
// ------------------------------------------------------------------------

// horizontal and vertical counters
reg [10:0]hcount;
reg [10:0]vcount;

// Horizontal and Vertical sync
reg HS,VS;

// active when inside visible screen area.
wire video_enable;

reg blank;


// increment horizontal counter at pixel_clk rate
// until HMAX is reached, then reset and keep counting
always @(posedge pixel_clk or negedge rst)
begin
 if(!rst)
  hcount <= 11'b0;
 else if(hcount == HMAX)
  hcount <= 11'b0;
 else
  hcount <= hcount + 1;
end

   
// increment vertical counter when one line is finished (horizontal counter reached HMAX)
// until VMAX is reached, then reset and keep counting
always @(posedge pixel_clk or negedge rst)
begin
 if(!rst)
  vcount <= 11'b0;
 else if(hcount == HMAX)
  begin
   if(vcount == VMAX)
    vcount <= 11'b0;
   else
    vcount <= vcount + 1;
  end
end


// generate horizontal synch pulse when horizontal counter is between where the
// front porch ends and the synch pulse ends.
// The HS is active (with polarity SPP) for a total of 96 pixels.
always @(posedge pixel_clk)
 begin
  if((hcount >= HFP) && (hcount < HSP))
    HS <= SPP;
  else
    HS <= !(SPP);
 end
  
	   
// generate vertical synch pulse when vertical counter is between where the
// front porch ends and the synch pulse ends.
// The VS is active (with polarity SPP) for a total of 2 video lines = 2*HMAX = 1600 pixels.
always @(posedge pixel_clk)
 begin
  if((vcount >= VFP) && (vcount < VSP))
    VS <= SPP;
  else
    VS <= !(SPP);
 end


// enable video output when pixel is in visible area
assign video_enable  = ((hcount < HLINES) && (vcount < VLINES)) ? 1'b1 : 1'b0;


// blank is active when outside screen visible area color output should be blacked (put on 0)
// when blank in active blank is delayed one pixel clock period from the video_enable
// signal to account for the pixel pipeline delay.
always @(posedge pixel_clk)
 blank <= !(video_enable);
 
     
endmodule
