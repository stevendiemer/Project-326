`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:10:47 03/08/2012 
// Design Name: 
// Module Name:    coin_driver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module coin_driver(
    input [9:0] player_left,
    input [9:0] player_right,
    output [3:0] coin_out
    );


endmodule
